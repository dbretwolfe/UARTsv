module Timing_Gen #(parameter SYSCLK_RATE = 100000000,
		parameter BAUD_RATE = 9600)
		
		(input logic SysClk,
		input Rst,
		output logic Clk);

	localparam CLOCK_DIV = SYSCLK_RATE / BAUD_RATE; // Baud rate is transitions per second.  We get one transition per rising
								// clock edge, meaning we need two clock transitions per baud.
	integer ClockCounter;

	always @ (posedge SysClk) begin
		if (ClockCounter === CLOCK_DIV - 1) begin
			Clk = ~Clk;
			ClockCounter = '0;
		end
		else begin
			Clk = Clk;
			ClockCounter = ClockCounter + 1;
		end
	end

endmodule