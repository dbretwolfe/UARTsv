module RX_FSM(Rx_In, Clk, Rst, RTS, Data_Rdy_Out, Rx_Data_Out, Rx_Error); 

parameter DATA_BITS = 9; // 8 data bits and one parity bit 
parameter STOP_BITS = 2;
parameter PARITY_BIT = 1;

input Rx_In;
input Clk;
input Rst;
output logic RTS;
output logic Data_Rdy_Out;
output logic [DATA_BITS-1:0] Rx_Data_Out;
output logic [2:0] Rx_Error;

logic [DATA_BITS-2:0] Data_Reg = 0; 
logic Parity_Bit=0;
logic [STOP_BITS-1:0] Reg_Stop = 0;
logic Reg_Parity =0;

int Count;
int Stop_Count;

enum {Ready, Start_Bit, Rx_Wait, Parity, Stop_Bit, Rx_Done } State, Next_State ; 	

always_ff @(posedge Clk)
begin 
	if(Rst) 
	State <= Ready;
	else 
	State <= Next_State;
end

always_comb
begin : set_Next_State

case(State)
	Ready: 	if(Rx_In == 0)
			Next_State =  Start_Bit;
		else
			Next_State = Ready;
	Start_Bit:
			Next_State =  Rx_Wait;
			
	Rx_Wait: 
		if (Count == DATA_BITS-1)
			Next_State = Parity;
		else 	
			Next_State = Rx_Wait;
			
	Parity  : 
			Next_State = Stop_Bit;
  	 
	Stop_Bit: 
		if(Stop_Count < STOP_BITS)
			Next_State = Stop_Bit;	
		else 
			Next_State = Rx_Done;
	Rx_Done: 	
		if(Rx_In == 1)
			Next_State = Ready;
		else
			Next_State = Rx_Done;
endcase;
end : set_Next_State;

always_comb
begin: set_Outputs	

	RTS = 1'b0;
	Rx_Error[2] = 1'b0;
	Rx_Error[1] = 1'b0;
	Rx_Error[0] = 1'b0;
	Rx_Data_Out = 0;
	Data_Rdy_Out = 0;

case(State)
	Ready: 
		 	RTS = 1'b1;
			
	Rx_Done: 	begin
			// Break Error 
			if((Data_Reg == 0) & (Reg_Stop != '1)) Rx_Error[0] = 1'b1;
			
			// Parity Error 
			for (int i = 1; i<DATA_BITS-1; i++)
				begin Parity_Bit = Data_Reg[i] ^ Data_Reg[i-1]; end
					if(Parity_Bit != Reg_Parity) Rx_Error[1] = 1'b1;
			
			// Framing Error 
			if(Reg_Stop != '1) Rx_Error[2] = 1'b1;
			
			// Data bits Output if there is no error in the data sent 
			if ( (Rx_Error[2] == 1'b1) | (Rx_Error[1] == 1'b1) |(Rx_Error[0] == 1'b1) )
				Rx_Data_Out = 0;
			else
				begin
				Rx_Data_Out = Data_Reg;		
				Data_Rdy_Out = 1;
				end
			end
endcase;
end : set_Outputs
 

always_ff @(posedge Clk)
begin 
if (Next_State == Ready ) 
begin
	Count = 0;
	Stop_Count=0;
	Data_Reg =0 ;
end
else if((Next_State == Rx_Wait) && (Count < DATA_BITS))
begin   
	Count = Count+1;
	Data_Reg = (Data_Reg << 1);
	Data_Reg = Data_Reg | Rx_In; 
end
else if (Next_State == Stop_Bit)
	begin
	Stop_Count = Stop_Count+1;
	Reg_Stop = (Reg_Stop <<1);
	Reg_Stop = Reg_Stop |Rx_In;
	end
else if (Next_State == Parity)
	Reg_Parity = Rx_In;
end
endmodule